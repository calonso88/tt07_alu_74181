module alu_74181_arith (a, b, s, f);

  input logic [3:0] a, b, s;
  output logic [3:0] f;

endmodule
